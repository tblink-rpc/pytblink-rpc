/*****************************************************************************
 * tblink.sv
 * TbLink SystemVerilog package
 *****************************************************************************/
package tblink;
	
	
	
endpackage
